module mutiplexGateLevel(A, B, X, out1);

input A, B, X;
output out1;

endmodule 
